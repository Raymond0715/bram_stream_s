`define WE_192			192'hffffffffffffffffffffffffffffffffffffffffffffffff
